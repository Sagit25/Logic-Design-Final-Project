`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:08:52 05/30/2022 
// Design Name: 
// Module Name:    hex7Segment 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module hex7Segment(
    input [7:0] input8Bit,
    output [13:0] LCDOutput
    );
	 
	 case(input8Bit) 
	 
	 endcase
	 


endmodule
